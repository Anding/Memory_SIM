library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


architecture sim of blk_mem_sim is

begin

end architecture;

